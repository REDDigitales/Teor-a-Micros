`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/18/2017 03:36:45 PM
// Design Name: 
// Module Name: Memoria_Principal
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Memoria_Principal(
    input clk,
    input Enable,
   EnMem,
   Dir_Instru,
   Dir_Mem,
   Dato_Instru,
   Dato_Mem
  
    );
endmodule
